class ncsu_void;

  function new(string name = ""); 
  endfunction

endclass
