virtual class ncsu_object_wrapper;
  pure virtual function string get_type_name();
  pure virtual function ncsu_object create_object(string name);
endclass
