package my_pkg;
	import ncsu_pkg::*;
	`include "ncsu_macros.svh"

	`include "src/transaction_handler.svh"
endpackage
